* c:\esim\fossee\esim\examples\jktod\jktod.cir

.lib "skywater-pdk-libs-sky130_fd_pr-main/models/sky130.lib.spice" tt
.include 3_and.sub
.include PMOS-0.5um.lib
.include NMOS-0.5um.lib
x1 net-_u1-pad3_ net-_u6-pad2_ net-_u1-pad4_ net-_u4-pad1_ 3_and
x2 net-_u1-pad4_ net-_u11-pad2_ net-_u6-pad3_ net-_u5-pad1_ 3_and
* u4  net-_u4-pad1_ net-_u4-pad2_ d_inverter
* u5  net-_u5-pad1_ net-_u5-pad2_ d_inverter
* u6  net-_u4-pad2_ net-_u6-pad2_ net-_u6-pad3_ d_nand
* u7  net-_u6-pad3_ net-_u5-pad2_ net-_u6-pad2_ d_nand
m2 net-_m1-pad1_ din vdd vdd sky130_fd_pr__pfet_01v8 W = 1.26, L = 0.15
m1 net-_m1-pad1_ din gnd gnd sky130_fd_pr__nfet_01v8 W = 1.26, L = 0.15
* u1  din clk net-_u1-pad3_ net-_u1-pad4_ adc_bridge_2
* u8  net-_u6-pad3_ net-_u6-pad2_ qout qnout dac_bridge_2
r2  qout gnd mid 1k sky130_fd_pr__res_generic_pd l=10
r1  qnout gnd mid 1k sky130_fd_pr__res_generic_pd l=10
v2  clk gnd pulse(0 5 1m 1m 1m 20 40)
* u10  qout plot_v1
* u9  qnout plot_v1
* u11  net-_m1-pad1_ net-_u11-pad2_ adc_bridge_1
* u2  din plot_v1
* u3  clk plot_v1
v1  vdd gnd 5
v3  din gnd pulse(0 5 1m 1m 1m 50 100)
a1 net-_u4-pad1_ net-_u4-pad2_ u4
a2 net-_u5-pad1_ net-_u5-pad2_ u5
a3 [net-_u4-pad2_ net-_u6-pad2_ ] net-_u6-pad3_ u6
a4 [net-_u6-pad3_ net-_u5-pad2_ ] net-_u6-pad2_ u7
a5 [din clk ] [net-_u1-pad3_ net-_u1-pad4_ ] u1
a6 [net-_u6-pad3_ net-_u6-pad2_ ] [qout qnout ] u8
a7 [net-_m1-pad1_ ] [net-_u11-pad2_ ] u11
* Schematic Name:                             d_inverter, NgSpice Name: d_inverter
.model u4 d_inverter(rise_delay=1.0e-9 fall_delay=1.0e-9 input_load=1.0e-12 ) 
* Schematic Name:                             d_inverter, NgSpice Name: d_inverter
.model u5 d_inverter(rise_delay=1.0e-9 fall_delay=1.0e-9 input_load=1.0e-12 ) 
* Schematic Name:                             d_nand, NgSpice Name: d_nand
.model u6 d_nand(rise_delay=1.0e-9 fall_delay=1.0e-9 input_load=1.0e-12 ) 
* Schematic Name:                             d_nand, NgSpice Name: d_nand
.model u7 d_nand(rise_delay=1.0e-9 fall_delay=1.0e-9 input_load=1.0e-12 ) 
* Schematic Name:                             adc_bridge_2, NgSpice Name: adc_bridge
.model u1 adc_bridge(in_low=1.0 in_high=2.0 rise_delay=1.0e-9 fall_delay=1.0e-9 ) 
* Schematic Name:                             dac_bridge_2, NgSpice Name: dac_bridge
.model u8 dac_bridge(out_low=0.0 out_high=5.0 out_undef=0.5 input_load=1.0e-12 t_rise=1.0e-9 t_fall=1.0e-9 ) 
* Schematic Name:                             adc_bridge_1, NgSpice Name: adc_bridge
.model u11 adc_bridge(in_low=1.0 in_high=2.0 rise_delay=1.0e-9 fall_delay=1.0e-9 ) 
.tran 10e-00 100e-00 0e-00

* Control Statements 
.control
run
print allv > plot_data_v.txt
print alli > plot_data_i.txt
plot v(qout)
plot v(qnout)
plot v(din)
plot v(clk)
.endc
.end
